VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM8
  CLASS BLOCK ;
  FOREIGN RAM8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 395.140 BY 27.200 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.140 4.120 395.140 4.720 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.140 6.840 395.140 7.440 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.140 9.560 395.140 10.160 ;
    END
  END A0[2]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.140 12.280 395.140 12.880 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 25.200 12.330 27.200 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 25.200 131.930 27.200 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 25.200 143.890 27.200 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 25.200 155.850 27.200 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 25.200 167.810 27.200 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 25.200 179.770 27.200 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 25.200 191.730 27.200 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 25.200 203.690 27.200 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 25.200 215.650 27.200 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 25.200 227.610 27.200 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 25.200 239.570 27.200 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 25.200 24.290 27.200 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 25.200 251.530 27.200 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 25.200 263.490 27.200 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 25.200 275.450 27.200 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 25.200 287.410 27.200 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 25.200 299.370 27.200 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 25.200 311.330 27.200 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 25.200 323.290 27.200 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 25.200 335.250 27.200 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 25.200 347.210 27.200 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 25.200 359.170 27.200 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 25.200 36.250 27.200 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 25.200 371.130 27.200 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 25.200 383.090 27.200 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 25.200 48.210 27.200 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 25.200 60.170 27.200 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 25.200 72.130 27.200 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 25.200 84.090 27.200 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 25.200 96.050 27.200 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 25.200 108.010 27.200 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 25.200 119.970 27.200 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.140 1.400 395.140 2.000 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 24.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 24.720 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 24.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 24.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 24.720 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.140 15.000 395.140 15.600 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.140 17.720 395.140 18.320 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.140 20.440 395.140 21.040 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 393.140 23.160 395.140 23.760 ;
    END
  END WE0[3]
  OBS
      LAYER nwell ;
        RECT 2.570 23.125 85.175 23.175 ;
        RECT 2.570 20.395 392.570 23.125 ;
        RECT 2.570 20.345 84.715 20.395 ;
        RECT 2.570 17.685 85.175 17.735 ;
        RECT 2.570 14.955 392.570 17.685 ;
        RECT 2.570 14.905 84.715 14.955 ;
        RECT 2.570 12.245 85.175 12.295 ;
        RECT 2.570 9.515 392.570 12.245 ;
        RECT 2.570 9.465 84.715 9.515 ;
        RECT 2.570 6.805 85.175 6.855 ;
        RECT 2.570 4.075 392.570 6.805 ;
        RECT 2.570 4.025 84.715 4.075 ;
      LAYER li1 ;
        RECT 2.760 2.635 392.380 24.565 ;
      LAYER met1 ;
        RECT 2.760 0.040 392.770 26.140 ;
      LAYER met2 ;
        RECT 4.700 24.920 11.770 26.170 ;
        RECT 12.610 24.920 23.730 26.170 ;
        RECT 24.570 24.920 35.690 26.170 ;
        RECT 36.530 24.920 47.650 26.170 ;
        RECT 48.490 24.920 59.610 26.170 ;
        RECT 60.450 24.920 71.570 26.170 ;
        RECT 72.410 24.920 83.530 26.170 ;
        RECT 84.370 24.920 95.490 26.170 ;
        RECT 96.330 24.920 107.450 26.170 ;
        RECT 108.290 24.920 119.410 26.170 ;
        RECT 120.250 24.920 131.370 26.170 ;
        RECT 132.210 24.920 143.330 26.170 ;
        RECT 144.170 24.920 155.290 26.170 ;
        RECT 156.130 24.920 167.250 26.170 ;
        RECT 168.090 24.920 179.210 26.170 ;
        RECT 180.050 24.920 191.170 26.170 ;
        RECT 192.010 24.920 203.130 26.170 ;
        RECT 203.970 24.920 215.090 26.170 ;
        RECT 215.930 24.920 227.050 26.170 ;
        RECT 227.890 24.920 239.010 26.170 ;
        RECT 239.850 24.920 250.970 26.170 ;
        RECT 251.810 24.920 262.930 26.170 ;
        RECT 263.770 24.920 274.890 26.170 ;
        RECT 275.730 24.920 286.850 26.170 ;
        RECT 287.690 24.920 298.810 26.170 ;
        RECT 299.650 24.920 310.770 26.170 ;
        RECT 311.610 24.920 322.730 26.170 ;
        RECT 323.570 24.920 334.690 26.170 ;
        RECT 335.530 24.920 346.650 26.170 ;
        RECT 347.490 24.920 358.610 26.170 ;
        RECT 359.450 24.920 370.570 26.170 ;
        RECT 371.410 24.920 382.530 26.170 ;
        RECT 383.370 24.920 392.750 26.170 ;
        RECT 4.700 2.280 392.750 24.920 ;
        RECT 4.700 0.010 11.770 2.280 ;
        RECT 12.610 0.010 23.730 2.280 ;
        RECT 24.570 0.010 35.690 2.280 ;
        RECT 36.530 0.010 47.650 2.280 ;
        RECT 48.490 0.010 59.610 2.280 ;
        RECT 60.450 0.010 71.570 2.280 ;
        RECT 72.410 0.010 83.530 2.280 ;
        RECT 84.370 0.010 95.490 2.280 ;
        RECT 96.330 0.010 107.450 2.280 ;
        RECT 108.290 0.010 119.410 2.280 ;
        RECT 120.250 0.010 131.370 2.280 ;
        RECT 132.210 0.010 143.330 2.280 ;
        RECT 144.170 0.010 155.290 2.280 ;
        RECT 156.130 0.010 167.250 2.280 ;
        RECT 168.090 0.010 179.210 2.280 ;
        RECT 180.050 0.010 191.170 2.280 ;
        RECT 192.010 0.010 203.130 2.280 ;
        RECT 203.970 0.010 215.090 2.280 ;
        RECT 215.930 0.010 227.050 2.280 ;
        RECT 227.890 0.010 239.010 2.280 ;
        RECT 239.850 0.010 250.970 2.280 ;
        RECT 251.810 0.010 262.930 2.280 ;
        RECT 263.770 0.010 274.890 2.280 ;
        RECT 275.730 0.010 286.850 2.280 ;
        RECT 287.690 0.010 298.810 2.280 ;
        RECT 299.650 0.010 310.770 2.280 ;
        RECT 311.610 0.010 322.730 2.280 ;
        RECT 323.570 0.010 334.690 2.280 ;
        RECT 335.530 0.010 346.650 2.280 ;
        RECT 347.490 0.010 358.610 2.280 ;
        RECT 359.450 0.010 370.570 2.280 ;
        RECT 371.410 0.010 382.530 2.280 ;
        RECT 383.370 0.010 392.750 2.280 ;
      LAYER met3 ;
        RECT 18.290 24.160 393.140 24.645 ;
        RECT 18.290 22.760 392.740 24.160 ;
        RECT 18.290 21.440 393.140 22.760 ;
        RECT 18.290 20.040 392.740 21.440 ;
        RECT 18.290 18.720 393.140 20.040 ;
        RECT 18.290 17.320 392.740 18.720 ;
        RECT 18.290 16.000 393.140 17.320 ;
        RECT 18.290 14.600 392.740 16.000 ;
        RECT 18.290 13.280 393.140 14.600 ;
        RECT 18.290 11.880 392.740 13.280 ;
        RECT 18.290 10.560 393.140 11.880 ;
        RECT 18.290 9.160 392.740 10.560 ;
        RECT 18.290 7.840 393.140 9.160 ;
        RECT 18.290 6.440 392.740 7.840 ;
        RECT 18.290 5.120 393.140 6.440 ;
        RECT 18.290 3.720 392.740 5.120 ;
        RECT 18.290 2.400 393.140 3.720 ;
        RECT 18.290 1.000 392.740 2.400 ;
        RECT 18.290 0.175 393.140 1.000 ;
      LAYER met4 ;
        RECT 282.735 4.935 325.080 20.905 ;
        RECT 327.480 4.935 375.065 20.905 ;
  END
END RAM8
END LIBRARY

